module vga_seven_segment (
    input clk,
    input [9:0] x,              // Current VGA x position
    input [9:0] y,              // Current VGA y position
    input [6:0] seg7_dig0,           // Rightmost digit (HEX0)
    input [6:0] seg7_dig1,           // HEX1
    input [6:0] seg7_dig2,           // HEX2
    input [6:0] seg7_dig3,           // HEX3
    input [6:0] seg7_dig4,           // Leftmost digit (HEX4)
    input [6:0] seg7_neg_sign,        // Negative sign (HEX5)
    output reg in_digit,             // High when pixel is part of a segment
    output reg [23:0] digit_color    // Color for the segment
);

// Display parameters
parameter BASE_X = 10'd10;       // Starting X position
parameter BASE_Y = 10'd405;      // Starting Y position
parameter DIGIT_WIDTH = 10'd30;  // Width of each digit
parameter DIGIT_HEIGHT = 10'd40; // Height of each digit
parameter DIGIT_SPACING = 10'd35; // Space between digits
parameter SEGMENT_THICKNESS = 10'd4; // Thickness of segments

// Segment colors
parameter SEG_ON_COLOR = 24'h000000;   // Red when on
parameter SEG_OFF_COLOR = 24'h006080;  // blue background when off

// Calculate which digit we're in
wire [9:0] digit_x [0:5];  // X position for each digit
assign digit_x[5] = BASE_X;
assign digit_x[4] = BASE_X + DIGIT_SPACING;
assign digit_x[3] = BASE_X + DIGIT_SPACING * 2;
assign digit_x[2] = BASE_X + DIGIT_SPACING * 3;
assign digit_x[1] = BASE_X + DIGIT_SPACING * 4;
assign digit_x[0] = BASE_X + DIGIT_SPACING * 5;

// Relative position within a digit
wire [9:0] rel_x;
wire [9:0] rel_y;
reg [2:0] current_digit;

// Seven segment layout (active low, so 0 = on)
// Segment positions:
//     aaa
//    f   b
//     ggg
//    e   c
//     ddd

wire [6:0] current_seg;
reg seg_a, seg_b, seg_c, seg_d, seg_e, seg_f, seg_g;

always @(*) begin
    in_digit = 0;
    current_digit = 3'd0;
    
    // Determine which digit position we're in
    if (y >= BASE_Y && y < BASE_Y + DIGIT_HEIGHT) begin
        if (x >= digit_x[5] && x < digit_x[5] + DIGIT_WIDTH) begin
            current_digit = 3'd5;
            in_digit = 1;
        end else if (x >= digit_x[4] && x < digit_x[4] + DIGIT_WIDTH) begin
            current_digit = 3'd4;
            in_digit = 1;
        end else if (x >= digit_x[3] && x < digit_x[3] + DIGIT_WIDTH) begin
            current_digit = 3'd3;
            in_digit = 1;
        end else if (x >= digit_x[2] && x < digit_x[2] + DIGIT_WIDTH) begin
            current_digit = 3'd2;
            in_digit = 1;
        end else if (x >= digit_x[1] && x < digit_x[1] + DIGIT_WIDTH) begin
            current_digit = 3'd1;
            in_digit = 1;
        end else if (x >= digit_x[0] && x < digit_x[0] + DIGIT_WIDTH) begin
            current_digit = 3'd0;
            in_digit = 1;
        end
    end
end

// Get relative coordinates within the digit
assign rel_x = x - digit_x[current_digit];
assign rel_y = y - BASE_Y;

// Select the appropriate segment data
assign current_seg = (current_digit == 3'd0) ? seg7_dig0 :
                     (current_digit == 3'd1) ? seg7_dig1 :
                     (current_digit == 3'd2) ? seg7_dig2 :
                     (current_digit == 3'd3) ? seg7_dig3 :
                     (current_digit == 3'd4) ? seg7_dig4 :
                     seg7_neg_sign;

// Extract individual segments (active low)
always @(*) begin
    seg_a = ~current_seg[0];
    seg_b = ~current_seg[1];
    seg_c = ~current_seg[2];
    seg_d = ~current_seg[3];
    seg_e = ~current_seg[4];
    seg_f = ~current_seg[5];
    seg_g = ~current_seg[6];
end

// Determine if current pixel is in any segment
reg in_seg_a, in_seg_b, in_seg_c, in_seg_d, in_seg_e, in_seg_f, in_seg_g;

always @(*) begin
    // Segment A (top horizontal)
    in_seg_a = (rel_y < SEGMENT_THICKNESS) && 
               (rel_x >= SEGMENT_THICKNESS) && 
               (rel_x < DIGIT_WIDTH - SEGMENT_THICKNESS);
    
    // Segment B (top right vertical)
    in_seg_b = (rel_y >= SEGMENT_THICKNESS) && 
               (rel_y < DIGIT_HEIGHT/2) &&
               (rel_x >= DIGIT_WIDTH - SEGMENT_THICKNESS);
    
    // Segment C (bottom right vertical)
    in_seg_c = (rel_y >= DIGIT_HEIGHT/2) && 
               (rel_y < DIGIT_HEIGHT - SEGMENT_THICKNESS) &&
               (rel_x >= DIGIT_WIDTH - SEGMENT_THICKNESS);
    
    // Segment D (bottom horizontal)
    in_seg_d = (rel_y >= DIGIT_HEIGHT - SEGMENT_THICKNESS) && 
               (rel_x >= SEGMENT_THICKNESS) && 
               (rel_x < DIGIT_WIDTH - SEGMENT_THICKNESS);
    
    // Segment E (bottom left vertical)
    in_seg_e = (rel_y >= DIGIT_HEIGHT/2) && 
               (rel_y < DIGIT_HEIGHT - SEGMENT_THICKNESS) &&
               (rel_x < SEGMENT_THICKNESS);
    
    // Segment F (top left vertical)
    in_seg_f = (rel_y >= SEGMENT_THICKNESS) && 
               (rel_y < DIGIT_HEIGHT/2) &&
               (rel_x < SEGMENT_THICKNESS);
    
    // Segment G (middle horizontal)
    in_seg_g = (rel_y >= DIGIT_HEIGHT/2 - SEGMENT_THICKNESS/2) && 
               (rel_y < DIGIT_HEIGHT/2 + SEGMENT_THICKNESS/2) &&
               (rel_x >= SEGMENT_THICKNESS) && 
               (rel_x < DIGIT_WIDTH - SEGMENT_THICKNESS);
    
    // Determine color based on which segment is active
    if (in_digit) begin
        if ((in_seg_a && seg_a) || (in_seg_b && seg_b) || 
            (in_seg_c && seg_c) || (in_seg_d && seg_d) ||
            (in_seg_e && seg_e) || (in_seg_f && seg_f) || 
            (in_seg_g && seg_g)) begin
            digit_color = SEG_ON_COLOR;
        end else if (in_seg_a || in_seg_b || in_seg_c || in_seg_d || 
                     in_seg_e || in_seg_f || in_seg_g) begin
            digit_color = SEG_OFF_COLOR;  // Show outline of off segments
        end else begin
            digit_color = 24'h006080;  // Background within digit area
        end
    end else begin
    digit_color = 24'h006080;
    end
end

endmodule