module timer(
input [9:0]timer,
output [6:0]timer_dig0,
output [6:0]timer_dig1,
output [6:0]timer_dig2
);

reg [3:0] result_one_digit;
reg [3:0] result_ten_digit;
reg [3:0] result_hundred_digit;

/* convert the binary value into 4 signals */
always @(*)
begin
		result_ten_digit = (timer / 10) % 10;
		result_one_digit = timer % 10;
		result_hundred_digit = (timer / 100) % 10;
end

/* instantiate the modules for each of the seven seg decoders including the negative one */
seven_segment dig2(.i(result_hundred_digit),.o(timer_dig2));
seven_segment dig1(.i(result_ten_digit),.o(timer_dig1));
seven_segment dig0(.i(result_one_digit),.o(timer_dig0));

endmodule